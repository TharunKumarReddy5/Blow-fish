`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:36:15 12/12/2013 
// Design Name: 
// Module Name:    s1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM( 
input[31:0] s1in,
input clk,rst,
output [31:0]sr1out
);
reg [31:0] s1out;
always @(s1in)
begin
case (s1in)
32'h00000000:s1out=32'hd1320ba6;
32'h00000001:s1out=32'h98dfb5ac;
32'h00000002:s1out=32'h2ffd72db;
32'h00000003:s1out=32'hd01adfb7;
32'h00000004:s1out=32'hb8e1afed;
32'h00000005:s1out=32'h6a267e96;
32'h00000006:s1out=32'hba7c9045;
32'h00000007:s1out=32'hf12c7f99;
32'h00000008:s1out=32'h24a19947;
32'h00000009:s1out=32'hb3916cf7;
32'h0000000a:s1out=32'h0801f2e2;
32'h0000000b:s1out=32'h858efc16;
32'h0000000c:s1out=32'h636920d8;
32'h0000000d:s1out=32'h71574e69;
32'h0000000e:s1out=32'ha458fea3;
32'h0000000f:s1out=32'hf4933d7e;

32'h00000010:s1out=32'h0d95748f;
32'h00000011:s1out=32'h728eb658;
32'h00000012:s1out=32'h718bcd58;
32'h00000013:s1out=32'h82154aee;
32'h00000014:s1out=32'h7b54a41d;
32'h00000015:s1out=32'hc25a59b5;
32'h00000016:s1out=32'h9c30d539;
32'h00000017:s1out=32'h2af26013;
32'h00000018:s1out=32'hc5d1b023;
32'h00000019:s1out=32'h286085f0;
32'h0000001a:s1out=32'hca417918;
32'h0000001b:s1out=32'hb8db38ef;
32'h0000001c:s1out=32'h8e79dcb0;
32'h0000001d:s1out=32'h603a180e;
32'h0000001e:s1out=32'h6c9e0e8b;
32'h0000001f:s1out=32'hb01e8a3e;

32'h00000020:s1out=32'hd71577c1;
32'h00000021:s1out=32'hbd324b27;
32'h00000022:s1out=32'h78af2fda;
32'h00000023:s1out=32'h55605c60;
32'h00000024:s1out=32'he65525f3;
32'h00000025:s1out=32'haa55ab94;
32'h00000026:s1out=32'h57489862;
32'h00000027:s1out=32'h63e81440;
32'h00000028:s1out=32'h55ca396a;
32'h00000029:s1out=32'h2aab10b6;
32'h0000002a:s1out=32'hb4cc5c34;
32'h0000002b:s1out=32'h1141e8ce;
32'h0000002c:s1out=32'ha15486af;
32'h0000002d:s1out=32'h7c72e993;
32'h0000002e:s1out=32'hb3ee1411;
32'h0000002f:s1out=32'h636fbc2a;

32'h00000030:s1out=32'h2ba9c55d;
32'h00000031:s1out=32'h741832f6;
32'h00000032:s1out=32'hce5c3e16;
32'h00000033:s1out=32'h9b87932e;
32'h00000034:s1out=32'hafd6ba33;
32'h00000035:s1out=32'h6c24cf5c;
32'h00000036:s1out=32'h7a325381;
32'h00000037:s1out=32'h28958677;
32'h00000038:s1out=32'h3b8f4898;
32'h00000039:s1out=32'h6b4bb9af;
32'h0000003a:s1out=32'hc4bfe81b;
32'h0000003b:s1out=32'h66282193;
32'h0000003c:s1out=32'h61d809cc;
32'h0000003d:s1out=32'hfb21a991;
32'h0000003e:s1out=32'h487cac60;
32'h0000003f:s1out=32'h5dec8032;

32'h00000040:s1out=32'hef845d5d;
32'h00000041:s1out=32'he98575b1;
32'h00000042:s1out=32'hdc262302;
32'h00000043:s1out=32'heb651b88;
32'h00000044:s1out=32'h23893e81;
32'h00000045:s1out=32'hd396acc5;
32'h00000046:s1out=32'h0f6d6ff3;
32'h00000047:s1out=32'h83f44239;
32'h00000048:s1out=32'h2e0b4482;
32'h00000049:s1out=32'ha4842004;
32'h0000004a:s1out=32'h69c8f04a;
32'h0000004b:s1out=32'h9e1f9b5e;
32'h0000004c:s1out=32'h21c66842;
32'h0000004d:s1out=32'hf6e96c9a;
32'h0000004e:s1out=32'h670c9c61;
32'h0000004f:s1out=32'habd388f0;

32'h00000050:s1out=32'h6a51a0d2;
32'h00000051:s1out=32'hd8542f68;
32'h00000052:s1out=32'h960fa728;
32'h00000053:s1out=32'hab5133a3;
32'h00000054:s1out=32'h6eef0b6c;
32'h00000055:s1out=32'h137a3be4;
32'h00000056:s1out=32'hba3bf050;
32'h00000057:s1out=32'h7efb2a98;
32'h00000058:s1out=32'ha1f1651d;
32'h00000059:s1out=32'h39af0176;
32'h0000005a:s1out=32'h66ca593e;
32'h0000005b:s1out=32'h82430e88;
32'h0000005c:s1out=32'h8cee8619;
32'h0000005d:s1out=32'h456f9fb4;
32'h0000005e:s1out=32'h7d84a5c3;
32'h0000005f:s1out=32'h3b8b5ebe;

32'h00000060:s1out=32'he06f75d8;
32'h00000061:s1out=32'h85c12073;
32'h00000062:s1out=32'h401a449f;
32'h00000063:s1out=32'h56c16aa6;
32'h00000064:s1out=32'h4ed3aa62;
32'h00000065:s1out=32'h363f7706;
32'h00000066:s1out=32'h1bfedf72;
32'h00000067:s1out=32'h429b023d;
32'h00000068:s1out=32'h37d0d724;
32'h00000069:s1out=32'hd00a1248;
32'h0000006a:s1out=32'hdb0fead3;
32'h0000006b:s1out=32'h49f1c09b;
32'h0000006c:s1out=32'h075372c9;
32'h0000006d:s1out=32'h80991b7b;
32'h0000006e:s1out=32'h25d479d8;
32'h0000006f:s1out=32'hf6e8def7;

32'h00000070:s1out=32'he3fe501a;
32'h00000071:s1out=32'hb6794c3b;
32'h00000072:s1out=32'h976ce0bd;
32'h00000073:s1out=32'h04c006ba;
32'h00000074:s1out=32'hc1a94fb6;
32'h00000075:s1out=32'h409f60c4;
32'h00000076:s1out=32'h5e5c9ec2;
32'h00000077:s1out=32'h196a2463;
32'h00000078:s1out=32'h68fb6faf;
32'h00000079:s1out=32'h3e6c53b5;
32'h0000007a:s1out=32'h1339b2eb;
32'h0000007b:s1out=32'h3b52ec6f;
32'h0000007c:s1out=32'h6dfc511f;
32'h0000007d:s1out=32'h9b30952c;
32'h0000007e:s1out=32'hcc814544;
32'h0000007f:s1out=32'haf5ebd09;

32'h00000080:s1out=32'hbee3d004;
32'h00000081:s1out=32'hde334afd;
32'h00000082:s1out=32'h660f2807;
32'h00000083:s1out=32'h192e4bb3;
32'h00000084:s1out=32'hc0cba857;
32'h00000085:s1out=32'h45c8740f;
32'h00000086:s1out=32'hd20b5f39;
32'h00000087:s1out=32'hb9d3fbdb;
32'h00000088:s1out=32'h5579c0bd;
32'h00000089:s1out=32'h1a60320a;
32'h0000008a:s1out=32'hd6a100c6;
32'h0000008b:s1out=32'h402c7279;
32'h0000008c:s1out=32'h679f25fe;
32'h0000008d:s1out=32'hfb1fa3cc;
32'h0000008e:s1out=32'h8ea5e9f8;
32'h0000008f:s1out=32'hdb3222f8;

32'h00000090:s1out=32'h3c7516df;
32'h00000091:s1out=32'hfd616b15;
32'h00000092:s1out=32'h2f501ec8;
32'h00000093:s1out=32'had0552ab;
32'h00000094:s1out=32'h323db5fa;
32'h00000095:s1out=32'hfd238760;
32'h00000096:s1out=32'h53327b48;
32'h00000097:s1out=32'h3e00df82;
32'h00000098:s1out=32'h9e5c57bb;
32'h00000099:s1out=32'hca6f8ca0;
32'h0000009a:s1out=32'h1a87562e;
32'h0000009b:s1out=32'hdf1769db;
32'h0000009c:s1out=32'hd542a8f6;
32'h0000009d:s1out=32'h287effc3;
32'h0000009e:s1out=32'hac6732c6;
32'h0000009f:s1out=32'h8c4f5573;

32'h000000a0:s1out=32'h695b27b0;
32'h000000a1:s1out=32'hbbca58c8;
32'h000000a2:s1out=32'he1ffa35d;
32'h000000a3:s1out=32'hb8f011a0;
32'h000000a4:s1out=32'h10fa3d98;
32'h000000a5:s1out=32'hfd2183b8;
32'h000000a6:s1out=32'h4afcb56c;
32'h000000a7:s1out=32'h2dd1d35b;
32'h000000a8:s1out=32'h9a53e479;
32'h000000a9:s1out=32'hb6f84565;
32'h000000aa:s1out=32'hd28e49bc;
32'h000000ab:s1out=32'h4bfb9790;
32'h000000ac:s1out=32'he1ddf2da;
32'h000000ad:s1out=32'ha4cb7e33;
32'h000000ae:s1out=32'h62fb1341;
32'h000000af:s1out=32'hcee4c6e8;

32'h000000b0:s1out=32'hef20cada;
32'h000000b1:s1out=32'h36774c01;
32'h000000b2:s1out=32'hd07e9efe;
32'h000000b3:s1out=32'h2bf11fb4;
32'h000000b4:s1out=32'h95dbda4d;
32'h000000b5:s1out=32'hae909198;
32'h000000b6:s1out=32'heaad8e71;
32'h000000b7:s1out=32'h6b93d5a0;
32'h000000b8:s1out=32'hd08ed1d0;
32'h000000b9:s1out=32'hafc725e0;
32'h000000ba:s1out=32'h8e3c5b2f;
32'h000000bb:s1out=32'h8e7594b7;
32'h000000bc:s1out=32'h8ff6e2fb;
32'h000000bd:s1out=32'hf2122b64;
32'h000000be:s1out=32'h8888b812;
32'h000000bf:s1out=32'h900df01c;

32'h000000c0:s1out=32'h4fad5ea0;
32'h000000c1:s1out=32'h688fc32c;
32'h000000c2:s1out=32'hd1cff191;
32'h000000c3:s1out=32'hb3a8c1ad;
32'h000000c4:s1out=32'h2f2f2218;
32'h000000c5:s1out=32'hbe0e1777;
32'h000000c6:s1out=32'hea752dfe;
32'h000000c7:s1out=32'h8b021fa1;
32'h000000c8:s1out=32'he5a0cc0f;
32'h000000c9:s1out=32'hb56f74e8;
32'h000000ca:s1out=32'h18acf3d6;
32'h000000cb:s1out=32'hce89e299;
32'h000000cc:s1out=32'hb4a84fe0;
32'h000000cd:s1out=32'hfd13e0b7;
32'h000000ce:s1out=32'h7cc43b81;
32'h000000cf:s1out=32'hd2ada8d9;

32'h000000d0:s1out=32'h165fa266;
32'h000000d1:s1out=32'h80957705;
32'h000000d2:s1out=32'h93cc7324;
32'h000000d3:s1out=32'h211a1477;
32'h000000d4:s1out=32'he6ad2065;
32'h000000d5:s1out=32'h77b5fa86;
32'h000000d6:s1out=32'hc75442f5;
32'h000000d7:s1out=32'hfb9d35cf;
32'h000000d8:s1out=32'hebcdaf0c;
32'h000000d9:s1out=32'h7b3e89a0;
32'h000000da:s1out=32'hd6411bd3;
32'h000000db:s1out=32'hae1e7e49;
32'h000000dc:s1out=32'h00250e2d;
32'h000000dd:s1out=32'h2071b35e;
32'h000000de:s1out=32'h226800bb;
32'h000000df:s1out=32'h57b8e0af;

32'h000000e0:s1out=32'h2464369b;
32'h000000e1:s1out=32'hf009b91e;
32'h000000e2:s1out=32'h5563911d;
32'h000000e3:s1out=32'h59dfa6aa;
32'h000000e4:s1out=32'h78c14389;
32'h000000e5:s1out=32'hd95a537f;
32'h000000e6:s1out=32'h207d5ba2;
32'h000000e7:s1out=32'h02e5b9c5;
32'h000000e8:s1out=32'h83260376;
32'h000000e9:s1out=32'h6295cfa9;
32'h000000ea:s1out=32'h11c81968;
32'h000000eb:s1out=32'h4e734a41;
32'h000000ec:s1out=32'hb3472dca;
32'h000000ed:s1out=32'h7b14a94a;
32'h000000ee:s1out=32'h1b510052;
32'h000000ef:s1out=32'h9a532915;

32'h000000f0:s1out=32'hd60f573f;
32'h000000f1:s1out=32'hbc9bc6e4;
32'h000000f2:s1out=32'h2b60a476;
32'h000000f3:s1out=32'h81e67400;
32'h000000f4:s1out=32'h08ba6fb5;
32'h000000f5:s1out=32'h571be91f;
32'h000000f6:s1out=32'hf296ec6b;
32'h000000f7:s1out=32'h2a0dd915;
32'h000000f8:s1out=32'hb6636521;
32'h000000f9:s1out=32'he7b9f9b6;
32'h000000fa:s1out=32'hff34052e;
32'h000000fb:s1out=32'hc5855664;
32'h000000fc:s1out=32'h53b02d5d;
32'h000000fd:s1out=32'ha99f8fa1;
32'h000000fe:s1out=32'h08ba4799;
32'h000000ff:s1out=32'h6e85076a;

//set2


32'h00000100:s1out=32'hd1320ba6;
32'h00000101:s1out=32'h98dfb5ac;
32'h00000102:s1out=32'h2ffd72db;
32'h00000103:s1out=32'hd01adfb7;
32'h00000104:s1out=32'hb8e1afed;
32'h00000105:s1out=32'h6a267e96;
32'h00000106:s1out=32'hba7c9045;
32'h00000107:s1out=32'hf12c7f99;
32'h00000108:s1out=32'h24a19947;
32'h00000109:s1out=32'hb3916cf7;
32'h0000010a:s1out=32'h0801f2e2;
32'h0000010b:s1out=32'h858efc16;
32'h0000010c:s1out=32'h636920d8;
32'h0000010d:s1out=32'h71574e69;
32'h0000010e:s1out=32'ha458fea3;
32'h0000010f:s1out=32'hf4933d7e;

32'h00000110:s1out=32'h0d95748f;
32'h00000111:s1out=32'h728eb658;
32'h00000112:s1out=32'h718bcd58;
32'h00000113:s1out=32'h82154aee;
32'h00000114:s1out=32'h7b54a41d;
32'h00000115:s1out=32'hc25a59b5;
32'h00000116:s1out=32'h9c30d539;
32'h00000117:s1out=32'h2af26013;
32'h00000118:s1out=32'hc5d1b023;
32'h00000119:s1out=32'h286085f0;
32'h0000011a:s1out=32'hca417918;
32'h0000011b:s1out=32'hb8db38ef;
32'h0000011c:s1out=32'h8e79dcb0;
32'h0000011d:s1out=32'h603a180e;
32'h0000011e:s1out=32'h6c9e0e8b;
32'h0000011f:s1out=32'hb01e8a3e;

32'h00000120:s1out=32'hd71577c1;
32'h00000121:s1out=32'hbd324b27;
32'h00000122:s1out=32'h78af2fda;
32'h00000123:s1out=32'h55605c60;
32'h00000124:s1out=32'he65525f3;
32'h00000125:s1out=32'haa55ab94;
32'h00000126:s1out=32'h57489862;
32'h00000127:s1out=32'h63e81440;
32'h00000128:s1out=32'h55ca396a;
32'h00000129:s1out=32'h2aab10b6;
32'h0000012a:s1out=32'hb4cc5c34;
32'h0000012b:s1out=32'h1141e8ce;
32'h0000012c:s1out=32'ha15486af;
32'h0000012d:s1out=32'h7c72e993;
32'h0000012e:s1out=32'hb3ee1411;
32'h0000012f:s1out=32'h636fbc2a;

32'h00000130:s1out=32'h2ba9c55d;
32'h00000131:s1out=32'h741832f6;
32'h00000132:s1out=32'hce5c3e16;
32'h00000133:s1out=32'h9b87932e;
32'h00000134:s1out=32'hafd6ba33;
32'h00000135:s1out=32'h6c24cf5c;
32'h00000136:s1out=32'h7a325381;
32'h00000137:s1out=32'h28958677;
32'h00000138:s1out=32'h3b8f4898;
32'h00000139:s1out=32'h6b4bb9af;
32'h0000013a:s1out=32'hc4bfe81b;
32'h0000013b:s1out=32'h66282193;
32'h0000013c:s1out=32'h61d809cc;
32'h0000013d:s1out=32'hfb21a991;
32'h0000013e:s1out=32'h487cac60;
32'h0000013f:s1out=32'h5dec8032;

32'h00000140:s1out=32'hef845d5d;
32'h00000141:s1out=32'he98575b1;
32'h00000142:s1out=32'hdc262302;
32'h00000143:s1out=32'heb651b88;
32'h00000144:s1out=32'h23893e81;
32'h00000145:s1out=32'hd396acc5;
32'h00000146:s1out=32'h0f6d6ff3;
32'h00000147:s1out=32'h83f44239;
32'h00000148:s1out=32'h2e0b4482;
32'h00000149:s1out=32'ha4842004;
32'h0000014a:s1out=32'h69c8f04a;
32'h0000014b:s1out=32'h9e1f9b5e;
32'h0000014c:s1out=32'h21c66842;
32'h0000014d:s1out=32'hf6e96c9a;
32'h0000014e:s1out=32'h670c9c61;
32'h0000014f:s1out=32'habd388f0;

32'h00000150:s1out=32'h6a51a0d2;
32'h00000151:s1out=32'hd8542f68;
32'h00000152:s1out=32'h960fa728;
32'h00000153:s1out=32'hab5133a3;
32'h00000154:s1out=32'h6eef0b6c;
32'h00000155:s1out=32'h137a3be4;
32'h00000156:s1out=32'hba3bf050;
32'h00000157:s1out=32'h7efb2a98;
32'h00000158:s1out=32'ha1f1651d;
32'h00000159:s1out=32'h39af0176;
32'h0000015a:s1out=32'h66ca593e;
32'h0000015b:s1out=32'h82430e88;
32'h0000015c:s1out=32'h8cee8619;
32'h0000015d:s1out=32'h456f9fb4;
32'h0000015e:s1out=32'h7d84a5c3;
32'h0000015f:s1out=32'h3b8b5ebe;

32'h00000160:s1out=32'he06f75d8;
32'h00000161:s1out=32'h85c12073;
32'h00000162:s1out=32'h401a449f;
32'h00000163:s1out=32'h56c16aa6;
32'h00000164:s1out=32'h4ed3aa62;
32'h00000165:s1out=32'h363f7706;
32'h00000166:s1out=32'h1bfedf72;
32'h00000167:s1out=32'h429b023d;
32'h00000168:s1out=32'h37d0d724;
32'h00000169:s1out=32'hd00a1248;
32'h0000016a:s1out=32'hdb0fead3;
32'h0000016b:s1out=32'h49f1c09b;
32'h0000016c:s1out=32'h075372c9;
32'h0000016d:s1out=32'h80991b7b;
32'h0000016e:s1out=32'h25d479d8;
32'h0000016f:s1out=32'hf6e8def7;

32'h00000170:s1out=32'he3fe501a;
32'h00000171:s1out=32'hb6794c3b;
32'h00000172:s1out=32'h976ce0bd;
32'h00000173:s1out=32'h04c006ba;
32'h00000174:s1out=32'hc1a94fb6;
32'h00000175:s1out=32'h409f60c4;
32'h00000176:s1out=32'h5e5c9ec2;
32'h00000177:s1out=32'h196a2463;
32'h00000178:s1out=32'h68fb6faf;
32'h00000179:s1out=32'h3e6c53b5;
32'h0000017a:s1out=32'h1339b2eb;
32'h0000017b:s1out=32'h3b52ec6f;
32'h0000017c:s1out=32'h6dfc511f;
32'h0000017d:s1out=32'h9b30952c;
32'h0000017e:s1out=32'hcc814544;
32'h0000017f:s1out=32'haf5ebd09;

32'h00000180:s1out=32'hbee3d004;
32'h00000181:s1out=32'hde334afd;
32'h00000182:s1out=32'h660f2807;
32'h00000183:s1out=32'h192e4bb3;
32'h00000184:s1out=32'hc0cba857;
32'h00000185:s1out=32'h45c8740f;
32'h00000186:s1out=32'hd20b5f39;
32'h00000187:s1out=32'hb9d3fbdb;
32'h00000188:s1out=32'h5579c0bd;
32'h00000189:s1out=32'h1a60320a;
32'h0000018a:s1out=32'hd6a100c6;
32'h0000018b:s1out=32'h402c7279;
32'h0000018c:s1out=32'h679f25fe;
32'h0000018d:s1out=32'hfb1fa3cc;
32'h0000018e:s1out=32'h8ea5e9f8;
32'h0000018f:s1out=32'hdb3222f8;

32'h00000190:s1out=32'h3c7516df;
32'h00000191:s1out=32'hfd616b15;
32'h00000192:s1out=32'h2f501ec8;
32'h00000193:s1out=32'had0552ab;
32'h00000194:s1out=32'h323db5fa;
32'h00000195:s1out=32'hfd238760;
32'h00000196:s1out=32'h53327b48;
32'h00000197:s1out=32'h3e00df82;
32'h00000198:s1out=32'h9e5c57bb;
32'h00000199:s1out=32'hca6f8ca0;
32'h0000019a:s1out=32'h1a87562e;
32'h0000019b:s1out=32'hdf1769db;
32'h0000019c:s1out=32'hd542a8f6;
32'h0000019d:s1out=32'h287effc3;
32'h0000019e:s1out=32'hac6732c6;
32'h0000019f:s1out=32'h8c4f5573;

32'h000001a0:s1out=32'h695b27b0;
32'h000001a1:s1out=32'hbbca58c8;
32'h000001a2:s1out=32'he1ffa35d;
32'h000001a3:s1out=32'hb8f011a0;
32'h000001a4:s1out=32'h10fa3d98;
32'h000001a5:s1out=32'hfd2183b8;
32'h000001a6:s1out=32'h4afcb56c;
32'h000001a7:s1out=32'h2dd1d35b;
32'h000001a8:s1out=32'h9a53e479;
32'h000001a9:s1out=32'hb6f84565;
32'h000001aa:s1out=32'hd28e49bc;
32'h000001ab:s1out=32'h4bfb9790;
32'h000001ac:s1out=32'he1ddf2da;
32'h000001ad:s1out=32'ha4cb7e33;
32'h000001ae:s1out=32'h62fb1341;
32'h000001af:s1out=32'hcee4c6e8;

32'h000001b0:s1out=32'hef20cada;
32'h000001b1:s1out=32'h36774c01;
32'h000001b2:s1out=32'hd07e9efe;
32'h000001b3:s1out=32'h2bf11fb4;
32'h000001b4:s1out=32'h95dbda4d;
32'h000001b5:s1out=32'hae909198;
32'h000001b6:s1out=32'heaad8e71;
32'h000001b7:s1out=32'h6b93d5a0;
32'h000001b8:s1out=32'hd08ed1d0;
32'h000001b9:s1out=32'hafc725e0;
32'h000001ba:s1out=32'h8e3c5b2f;
32'h000001bb:s1out=32'h8e7594b7;
32'h000001bc:s1out=32'h8ff6e2fb;
32'h000001bd:s1out=32'hf2122b64;
32'h000001be:s1out=32'h8888b812;
32'h000001bf:s1out=32'h900df01c;

32'h000001c0:s1out=32'h4fad5ea0;
32'h000001c1:s1out=32'h688fc32c;
32'h000001c2:s1out=32'hd1cff191;
32'h000001c3:s1out=32'hb3a8c1ad;
32'h000001c4:s1out=32'h2f2f2218;
32'h000001c5:s1out=32'hbe0e1777;
32'h000001c6:s1out=32'hea752dfe;
32'h000001c7:s1out=32'h8b021fa1;
32'h000001c8:s1out=32'he5a0cc0f;
32'h000001c9:s1out=32'hb56f74e8;
32'h000001ca:s1out=32'h18acf3d6;
32'h000001cb:s1out=32'hce89e299;
32'h000001cc:s1out=32'hb4a84fe0;
32'h000001cd:s1out=32'hfd13e0b7;
32'h000001ce:s1out=32'h7cc43b81;
32'h000001cf:s1out=32'hd2ada8d9;

32'h000001d0:s1out=32'h165fa266;
32'h000001d1:s1out=32'h80957705;
32'h000001d2:s1out=32'h93cc7324;
32'h000001d3:s1out=32'h211a1477;
32'h000001d4:s1out=32'he6ad2065;
32'h000001d5:s1out=32'h77b5fa86;
32'h000001d6:s1out=32'hc75442f5;
32'h000001d7:s1out=32'hfb9d35cf;
32'h000001d8:s1out=32'hebcdaf0c;
32'h000001d9:s1out=32'h7b3e89a0;
32'h000001da:s1out=32'hd6411bd3;
32'h000001db:s1out=32'hae1e7e49;
32'h000001dc:s1out=32'h00250e2d;
32'h000001dd:s1out=32'h2071b35e;
32'h000001de:s1out=32'h226800bb;
32'h000001df:s1out=32'h57b8e0af;

32'h000001e0:s1out=32'h2464369b;
32'h000001e1:s1out=32'hf009b91e;
32'h000001e2:s1out=32'h5563911d;
32'h000001e3:s1out=32'h59dfa6aa;
32'h000001e4:s1out=32'h78c14389;
32'h000001e5:s1out=32'hd95a537f;
32'h000001e6:s1out=32'h207d5ba2;
32'h000001e7:s1out=32'h02e5b9c5;
32'h000001e8:s1out=32'h83260376;
32'h000001e9:s1out=32'h6295cfa9;
32'h000001ea:s1out=32'h11c81968;
32'h000001eb:s1out=32'h4e734a41;
32'h000001ec:s1out=32'hb3472dca;
32'h000001ed:s1out=32'h7b14a94a;
32'h000001ee:s1out=32'h1b510052;
32'h000001ef:s1out=32'h9a532915;

32'h000001f0:s1out=32'hd60f573f;
32'h000001f1:s1out=32'hbc9bc6e4;
32'h000001f2:s1out=32'h2b60a476;
32'h000001f3:s1out=32'h81e67400;
32'h000001f4:s1out=32'h08ba6fb5;
32'h000001f5:s1out=32'h571be91f;
32'h000001f6:s1out=32'hf296ec6b;
32'h000001f7:s1out=32'h2a0dd915;
32'h000001f8:s1out=32'hb6636521;
32'h000001f9:s1out=32'he7b9f9b6;
32'h000001fa:s1out=32'hff34052e;
32'h000001fb:s1out=32'hc5855664;
32'h000001fc:s1out=32'h53b02d5d;
32'h000001fd:s1out=32'ha99f8fa1;
32'h000001fe:s1out=32'h08ba4799;
32'h000001ff:s1out=32'h6e85076a;

//set3


32'h00000200:s1out=32'hd1320ba6;
32'h00000201:s1out=32'h98dfb5ac;
32'h00000202:s1out=32'h2ffd72db;
32'h00000203:s1out=32'hd01adfb7;
32'h00000204:s1out=32'hb8e1afed;
32'h00000205:s1out=32'h6a267e96;
32'h00000206:s1out=32'hba7c9045;
32'h00000207:s1out=32'hf12c7f99;
32'h00000208:s1out=32'h24a19947;
32'h00000209:s1out=32'hb3916cf7;
32'h0000020a:s1out=32'h0801f2e2;
32'h0000020b:s1out=32'h858efc16;
32'h0000020c:s1out=32'h636920d8;
32'h0000020d:s1out=32'h71574e69;
32'h0000020e:s1out=32'ha458fea3;
32'h0000020f:s1out=32'hf4933d7e;

32'h00000210:s1out=32'h0d95748f;
32'h00000211:s1out=32'h728eb658;
32'h00000212:s1out=32'h718bcd58;
32'h00000213:s1out=32'h82154aee;
32'h00000214:s1out=32'h7b54a41d;
32'h00000215:s1out=32'hc25a59b5;
32'h00000216:s1out=32'h9c30d539;
32'h00000217:s1out=32'h2af26013;
32'h00000218:s1out=32'hc5d1b023;
32'h00000219:s1out=32'h286085f0;
32'h0000021a:s1out=32'hca417918;
32'h0000021b:s1out=32'hb8db38ef;
32'h0000021c:s1out=32'h8e79dcb0;
32'h0000021d:s1out=32'h603a180e;
32'h0000021e:s1out=32'h6c9e0e8b;
32'h0000021f:s1out=32'hb01e8a3e;

32'h00000220:s1out=32'hd71577c1;
32'h00000221:s1out=32'hbd324b27;
32'h00000222:s1out=32'h78af2fda;
32'h00000223:s1out=32'h55605c60;
32'h00000224:s1out=32'he65525f3;
32'h00000225:s1out=32'haa55ab94;
32'h00000226:s1out=32'h57489862;
32'h00000227:s1out=32'h63e81440;
32'h00000228:s1out=32'h55ca396a;
32'h00000229:s1out=32'h2aab10b6;
32'h0000022a:s1out=32'hb4cc5c34;
32'h0000022b:s1out=32'h1141e8ce;
32'h0000022c:s1out=32'ha15486af;
32'h0000022d:s1out=32'h7c72e993;
32'h0000022e:s1out=32'hb3ee1411;
32'h0000022f:s1out=32'h636fbc2a;

32'h00000230:s1out=32'h2ba9c55d;
32'h00000231:s1out=32'h741832f6;
32'h00000232:s1out=32'hce5c3e16;
32'h00000233:s1out=32'h9b87932e;
32'h00000234:s1out=32'hafd6ba33;
32'h00000235:s1out=32'h6c24cf5c;
32'h00000236:s1out=32'h7a325381;
32'h00000237:s1out=32'h28958677;
32'h00000238:s1out=32'h3b8f4898;
32'h00000239:s1out=32'h6b4bb9af;
32'h0000023a:s1out=32'hc4bfe81b;
32'h0000023b:s1out=32'h66282193;
32'h0000023c:s1out=32'h61d809cc;
32'h0000023d:s1out=32'hfb21a991;
32'h0000023e:s1out=32'h487cac60;
32'h0000023f:s1out=32'h5dec8032;

32'h00000240:s1out=32'hef845d5d;
32'h00000241:s1out=32'he98575b1;
32'h00000242:s1out=32'hdc262302;
32'h00000243:s1out=32'heb651b88;
32'h00000244:s1out=32'h23893e81;
32'h00000245:s1out=32'hd396acc5;
32'h00000246:s1out=32'h0f6d6ff3;
32'h00000247:s1out=32'h83f44239;
32'h00000248:s1out=32'h2e0b4482;
32'h00000249:s1out=32'ha4842004;
32'h0000024a:s1out=32'h69c8f04a;
32'h0000024b:s1out=32'h9e1f9b5e;
32'h0000024c:s1out=32'h21c66842;
32'h0000024d:s1out=32'hf6e96c9a;
32'h0000024e:s1out=32'h670c9c61;
32'h0000024f:s1out=32'habd388f0;

32'h00000250:s1out=32'h6a51a0d2;
32'h00000251:s1out=32'hd8542f68;
32'h00000252:s1out=32'h960fa728;
32'h00000253:s1out=32'hab5133a3;
32'h00000254:s1out=32'h6eef0b6c;
32'h00000255:s1out=32'h137a3be4;
32'h00000256:s1out=32'hba3bf050;
32'h00000257:s1out=32'h7efb2a98;
32'h00000258:s1out=32'ha1f1651d;
32'h00000259:s1out=32'h39af0176;
32'h0000025a:s1out=32'h66ca593e;
32'h0000025b:s1out=32'h82430e88;
32'h0000025c:s1out=32'h8cee8619;
32'h0000025d:s1out=32'h456f9fb4;
32'h0000025e:s1out=32'h7d84a5c3;
32'h0000025f:s1out=32'h3b8b5ebe;

32'h00000260:s1out=32'he06f75d8;
32'h00000261:s1out=32'h85c12073;
32'h00000262:s1out=32'h401a449f;
32'h00000263:s1out=32'h56c16aa6;
32'h00000264:s1out=32'h4ed3aa62;
32'h00000265:s1out=32'h363f7706;
32'h00000266:s1out=32'h1bfedf72;
32'h00000267:s1out=32'h429b023d;
32'h00000268:s1out=32'h37d0d724;
32'h00000269:s1out=32'hd00a1248;
32'h0000026a:s1out=32'hdb0fead3;
32'h0000026b:s1out=32'h49f1c09b;
32'h0000026c:s1out=32'h075372c9;
32'h0000026d:s1out=32'h80991b7b;
32'h0000026e:s1out=32'h25d479d8;
32'h0000026f:s1out=32'hf6e8def7;

32'h00000270:s1out=32'he3fe501a;
32'h00000271:s1out=32'hb6794c3b;
32'h00000272:s1out=32'h976ce0bd;
32'h00000273:s1out=32'h04c006ba;
32'h00000274:s1out=32'hc1a94fb6;
32'h00000275:s1out=32'h409f60c4;
32'h00000276:s1out=32'h5e5c9ec2;
32'h00000277:s1out=32'h196a2463;
32'h00000278:s1out=32'h68fb6faf;
32'h00000279:s1out=32'h3e6c53b5;
32'h0000027a:s1out=32'h1339b2eb;
32'h0000027b:s1out=32'h3b52ec6f;
32'h0000027c:s1out=32'h6dfc511f;
32'h0000027d:s1out=32'h9b30952c;
32'h0000027e:s1out=32'hcc814544;
32'h0000027f:s1out=32'haf5ebd09;

32'h00000280:s1out=32'hbee3d004;
32'h00000281:s1out=32'hde334afd;
32'h00000282:s1out=32'h660f2807;
32'h00000283:s1out=32'h192e4bb3;
32'h00000284:s1out=32'hc0cba857;
32'h00000285:s1out=32'h45c8740f;
32'h00000286:s1out=32'hd20b5f39;
32'h00000287:s1out=32'hb9d3fbdb;
32'h00000288:s1out=32'h5579c0bd;
32'h00000289:s1out=32'h1a60320a;
32'h0000028a:s1out=32'hd6a100c6;
32'h0000028b:s1out=32'h402c7279;
32'h0000028c:s1out=32'h679f25fe;
32'h0000028d:s1out=32'hfb1fa3cc;
32'h0000028e:s1out=32'h8ea5e9f8;
32'h0000028f:s1out=32'hdb3222f8;

32'h00000290:s1out=32'h3c7516df;
32'h00000291:s1out=32'hfd616b15;
32'h00000292:s1out=32'h2f501ec8;
32'h00000293:s1out=32'had0552ab;
32'h00000294:s1out=32'h323db5fa;
32'h00000295:s1out=32'hfd238760;
32'h00000296:s1out=32'h53327b48;
32'h00000297:s1out=32'h3e00df82;
32'h00000298:s1out=32'h9e5c57bb;
32'h00000299:s1out=32'hca6f8ca0;
32'h0000029a:s1out=32'h1a87562e;
32'h0000029b:s1out=32'hdf1769db;
32'h0000029c:s1out=32'hd542a8f6;
32'h0000029d:s1out=32'h287effc3;
32'h0000029e:s1out=32'hac6732c6;
32'h0000029f:s1out=32'h8c4f5573;

32'h000002a0:s1out=32'h695b27b0;
32'h000002a1:s1out=32'hbbca58c8;
32'h000002a2:s1out=32'he1ffa35d;
32'h000002a3:s1out=32'hb8f011a0;
32'h000002a4:s1out=32'h10fa3d98;
32'h000002a5:s1out=32'hfd2183b8;
32'h000002a6:s1out=32'h4afcb56c;
32'h000002a7:s1out=32'h2dd1d35b;
32'h000002a8:s1out=32'h9a53e479;
32'h000002a9:s1out=32'hb6f84565;
32'h000002aa:s1out=32'hd28e49bc;
32'h000002ab:s1out=32'h4bfb9790;
32'h000002ac:s1out=32'he1ddf2da;
32'h000002ad:s1out=32'ha4cb7e33;
32'h000002ae:s1out=32'h62fb1341;
32'h000002af:s1out=32'hcee4c6e8;

32'h000002b0:s1out=32'hef20cada;
32'h000002b1:s1out=32'h36774c01;
32'h000002b2:s1out=32'hd07e9efe;
32'h000002b3:s1out=32'h2bf11fb4;
32'h000002b4:s1out=32'h95dbda4d;
32'h000002b5:s1out=32'hae909198;
32'h000002b6:s1out=32'heaad8e71;
32'h000002b7:s1out=32'h6b93d5a0;
32'h000002b8:s1out=32'hd08ed1d0;
32'h000002b9:s1out=32'hafc725e0;
32'h000002ba:s1out=32'h8e3c5b2f;
32'h000002bb:s1out=32'h8e7594b7;
32'h000002bc:s1out=32'h8ff6e2fb;
32'h000002bd:s1out=32'hf2122b64;
32'h000002be:s1out=32'h8888b812;
32'h000002bf:s1out=32'h900df01c;

32'h000002c0:s1out=32'h4fad5ea0;
32'h000002c1:s1out=32'h688fc32c;
32'h000002c2:s1out=32'hd1cff191;
32'h000002c3:s1out=32'hb3a8c1ad;
32'h000002c4:s1out=32'h2f2f2218;
32'h000002c5:s1out=32'hbe0e1777;
32'h000002c6:s1out=32'hea752dfe;
32'h000002c7:s1out=32'h8b021fa1;
32'h000002c8:s1out=32'he5a0cc0f;
32'h000002c9:s1out=32'hb56f74e8;
32'h000002ca:s1out=32'h18acf3d6;
32'h000002cb:s1out=32'hce89e299;
32'h000002cc:s1out=32'hb4a84fe0;
32'h000002cd:s1out=32'hfd13e0b7;
32'h000002ce:s1out=32'h7cc43b81;
32'h000002cf:s1out=32'hd2ada8d9;

32'h000002d0:s1out=32'h165fa266;
32'h000002d1:s1out=32'h80957705;
32'h000002d2:s1out=32'h93cc7324;
32'h000002d3:s1out=32'h211a1477;
32'h000002d4:s1out=32'he6ad2065;
32'h000002d5:s1out=32'h77b5fa86;
32'h000002d6:s1out=32'hc75442f5;
32'h000002d7:s1out=32'hfb9d35cf;
32'h000002d8:s1out=32'hebcdaf0c;
32'h000002d9:s1out=32'h7b3e89a0;
32'h000002da:s1out=32'hd6411bd3;
32'h000002db:s1out=32'hae1e7e49;
32'h000002dc:s1out=32'h00250e2d;
32'h000002dd:s1out=32'h2071b35e;
32'h000002de:s1out=32'h226800bb;
32'h000002df:s1out=32'h57b8e0af;

32'h000002e0:s1out=32'h2464369b;
32'h000002e1:s1out=32'hf009b91e;
32'h000002e2:s1out=32'h5563911d;
32'h000002e3:s1out=32'h59dfa6aa;
32'h000002e4:s1out=32'h78c14389;
32'h000002e5:s1out=32'hd95a537f;
32'h000002e6:s1out=32'h207d5ba2;
32'h000002e7:s1out=32'h02e5b9c5;
32'h000002e8:s1out=32'h83260376;
32'h000002e9:s1out=32'h6295cfa9;
32'h000002ea:s1out=32'h11c81968;
32'h000002eb:s1out=32'h4e734a41;
32'h000002ec:s1out=32'hb3472dca;
32'h000002ed:s1out=32'h7b14a94a;
32'h000002ee:s1out=32'h1b510052;
32'h000002ef:s1out=32'h9a532915;

32'h000002f0:s1out=32'hd60f573f;
32'h000002f1:s1out=32'hbc9bc6e4;
32'h000002f2:s1out=32'h2b60a476;
32'h000002f3:s1out=32'h81e67400;
32'h000002f4:s1out=32'h08ba6fb5;
32'h000002f5:s1out=32'h571be91f;
32'h000002f6:s1out=32'hf296ec6b;
32'h000002f7:s1out=32'h2a0dd915;
32'h000002f8:s1out=32'hb6636521;
32'h000002f9:s1out=32'he7b9f9b6;
32'h000002fa:s1out=32'hff34052e;
32'h000002fb:s1out=32'hc5855664;
32'h000002fc:s1out=32'h53b02d5d;
32'h000002fd:s1out=32'ha99f8fa1;
32'h000002fe:s1out=32'h08ba4799;
32'h000002ff:s1out=32'h6e85076a;

//set4


32'h00000300:s1out=32'hd1320ba6;
32'h00000301:s1out=32'h98dfb5ac;
32'h00000302:s1out=32'h2ffd72db;
32'h00000303:s1out=32'hd01adfb7;
32'h00000304:s1out=32'hb8e1afed;
32'h00000305:s1out=32'h6a267e96;
32'h00000306:s1out=32'hba7c9045;
32'h00000307:s1out=32'hf12c7f99;
32'h00000308:s1out=32'h24a19947;
32'h00000309:s1out=32'hb3916cf7;
32'h0000030a:s1out=32'h0801f2e2;
32'h0000030b:s1out=32'h858efc16;
32'h0000030c:s1out=32'h636920d8;
32'h0000030d:s1out=32'h71574e69;
32'h0000030e:s1out=32'ha458fea3;
32'h0000030f:s1out=32'hf4933d7e;

32'h00000310:s1out=32'h0d95748f;
32'h00000311:s1out=32'h728eb658;
32'h00000312:s1out=32'h718bcd58;
32'h00000313:s1out=32'h82154aee;
32'h00000314:s1out=32'h7b54a41d;
32'h00000315:s1out=32'hc25a59b5;
32'h00000316:s1out=32'h9c30d539;
32'h00000317:s1out=32'h2af26013;
32'h00000318:s1out=32'hc5d1b023;
32'h00000319:s1out=32'h286085f0;
32'h0000031a:s1out=32'hca417918;
32'h0000031b:s1out=32'hb8db38ef;
32'h0000031c:s1out=32'h8e79dcb0;
32'h0000031d:s1out=32'h603a180e;
32'h0000031e:s1out=32'h6c9e0e8b;
32'h0000031f:s1out=32'hb01e8a3e;

32'h00000320:s1out=32'hd71577c1;
32'h00000321:s1out=32'hbd324b27;
32'h00000322:s1out=32'h78af2fda;
32'h00000323:s1out=32'h55605c60;
32'h00000324:s1out=32'he65525f3;
32'h00000325:s1out=32'haa55ab94;
32'h00000326:s1out=32'h57489862;
32'h00000327:s1out=32'h63e81440;
32'h00000328:s1out=32'h55ca396a;
32'h00000329:s1out=32'h2aab10b6;
32'h0000032a:s1out=32'hb4cc5c34;
32'h0000032b:s1out=32'h1141e8ce;
32'h0000032c:s1out=32'ha15486af;
32'h0000032d:s1out=32'h7c72e993;
32'h0000032e:s1out=32'hb3ee1411;
32'h0000032f:s1out=32'h636fbc2a;

32'h00000330:s1out=32'h2ba9c55d;
32'h00000331:s1out=32'h741832f6;
32'h00000332:s1out=32'hce5c3e16;
32'h00000333:s1out=32'h9b87932e;
32'h00000334:s1out=32'hafd6ba33;
32'h00000335:s1out=32'h6c24cf5c;
32'h00000336:s1out=32'h7a325381;
32'h00000337:s1out=32'h28958677;
32'h00000338:s1out=32'h3b8f4898;
32'h00000339:s1out=32'h6b4bb9af;
32'h0000033a:s1out=32'hc4bfe81b;
32'h0000033b:s1out=32'h66282193;
32'h0000033c:s1out=32'h61d809cc;
32'h0000033d:s1out=32'hfb21a991;
32'h0000033e:s1out=32'h487cac60;
32'h0000033f:s1out=32'h5dec8032;

32'h00000340:s1out=32'hef845d5d;
32'h00000341:s1out=32'he98575b1;
32'h00000342:s1out=32'hdc262302;
32'h00000343:s1out=32'heb651b88;
32'h00000344:s1out=32'h23893e81;
32'h00000345:s1out=32'hd396acc5;
32'h00000346:s1out=32'h0f6d6ff3;
32'h00000347:s1out=32'h83f44239;
32'h00000348:s1out=32'h2e0b4482;
32'h00000349:s1out=32'ha4842004;
32'h0000034a:s1out=32'h69c8f04a;
32'h0000034b:s1out=32'h9e1f9b5e;
32'h0000034c:s1out=32'h21c66842;
32'h0000034d:s1out=32'hf6e96c9a;
32'h0000034e:s1out=32'h670c9c61;
32'h0000034f:s1out=32'habd388f0;

32'h00000350:s1out=32'h6a51a0d2;
32'h00000351:s1out=32'hd8542f68;
32'h00000352:s1out=32'h960fa728;
32'h00000353:s1out=32'hab5133a3;
32'h00000354:s1out=32'h6eef0b6c;
32'h00000355:s1out=32'h137a3be4;
32'h00000356:s1out=32'hba3bf050;
32'h00000357:s1out=32'h7efb2a98;
32'h00000358:s1out=32'ha1f1651d;
32'h00000359:s1out=32'h39af0176;
32'h0000035a:s1out=32'h66ca593e;
32'h0000035b:s1out=32'h82430e88;
32'h0000035c:s1out=32'h8cee8619;
32'h0000035d:s1out=32'h456f9fb4;
32'h0000035e:s1out=32'h7d84a5c3;
32'h0000035f:s1out=32'h3b8b5ebe;

32'h00000360:s1out=32'he06f75d8;
32'h00000361:s1out=32'h85c12073;
32'h00000362:s1out=32'h401a449f;
32'h00000363:s1out=32'h56c16aa6;
32'h00000364:s1out=32'h4ed3aa62;
32'h00000365:s1out=32'h363f7706;
32'h00000366:s1out=32'h1bfedf72;
32'h00000367:s1out=32'h429b023d;
32'h00000368:s1out=32'h37d0d724;
32'h00000369:s1out=32'hd00a1248;
32'h0000036a:s1out=32'hdb0fead3;
32'h0000036b:s1out=32'h49f1c09b;
32'h0000036c:s1out=32'h075372c9;
32'h0000036d:s1out=32'h80991b7b;
32'h0000036e:s1out=32'h25d479d8;
32'h0000036f:s1out=32'hf6e8def7;

32'h00000370:s1out=32'he3fe501a;
32'h00000371:s1out=32'hb6794c3b;
32'h00000372:s1out=32'h976ce0bd;
32'h00000373:s1out=32'h04c006ba;
32'h00000374:s1out=32'hc1a94fb6;
32'h00000375:s1out=32'h409f60c4;
32'h00000376:s1out=32'h5e5c9ec2;
32'h00000377:s1out=32'h196a2463;
32'h00000378:s1out=32'h68fb6faf;
32'h00000379:s1out=32'h3e6c53b5;
32'h0000037a:s1out=32'h1339b2eb;
32'h0000037b:s1out=32'h3b52ec6f;
32'h0000037c:s1out=32'h6dfc511f;
32'h0000037d:s1out=32'h9b30952c;
32'h0000037e:s1out=32'hcc814544;
32'h0000037f:s1out=32'haf5ebd09;

32'h00000380:s1out=32'hbee3d004;
32'h00000381:s1out=32'hde334afd;
32'h00000382:s1out=32'h660f2807;
32'h00000383:s1out=32'h192e4bb3;
32'h00000384:s1out=32'hc0cba857;
32'h00000385:s1out=32'h45c8740f;
32'h00000386:s1out=32'hd20b5f39;
32'h00000387:s1out=32'hb9d3fbdb;
32'h00000388:s1out=32'h5579c0bd;
32'h00000389:s1out=32'h1a60320a;
32'h0000038a:s1out=32'hd6a100c6;
32'h0000038b:s1out=32'h402c7279;
32'h0000038c:s1out=32'h679f25fe;
32'h0000038d:s1out=32'hfb1fa3cc;
32'h0000038e:s1out=32'h8ea5e9f8;
32'h0000038f:s1out=32'hdb3222f8;

32'h00000390:s1out=32'h3c7516df;
32'h00000391:s1out=32'hfd616b15;
32'h00000392:s1out=32'h2f501ec8;
32'h00000393:s1out=32'had0552ab;
32'h00000394:s1out=32'h323db5fa;
32'h00000395:s1out=32'hfd238760;
32'h00000396:s1out=32'h53327b48;
32'h00000397:s1out=32'h3e00df82;
32'h00000398:s1out=32'h9e5c57bb;
32'h00000399:s1out=32'hca6f8ca0;
32'h0000039a:s1out=32'h1a87562e;
32'h0000039b:s1out=32'hdf1769db;
32'h0000039c:s1out=32'hd542a8f6;
32'h0000039d:s1out=32'h287effc3;
32'h0000039e:s1out=32'hac6732c6;
32'h0000039f:s1out=32'h8c4f5573;

32'h000003a0:s1out=32'h695b27b0;
32'h000003a1:s1out=32'hbbca58c8;
32'h000003a2:s1out=32'he1ffa35d;
32'h000003a3:s1out=32'hb8f011a0;
32'h000003a4:s1out=32'h10fa3d98;
32'h000003a5:s1out=32'hfd2183b8;
32'h000003a6:s1out=32'h4afcb56c;
32'h000003a7:s1out=32'h2dd1d35b;
32'h000003a8:s1out=32'h9a53e479;
32'h000003a9:s1out=32'hb6f84565;
32'h000003aa:s1out=32'hd28e49bc;
32'h000003ab:s1out=32'h4bfb9790;
32'h000003ac:s1out=32'he1ddf2da;
32'h000003ad:s1out=32'ha4cb7e33;
32'h000003ae:s1out=32'h62fb1341;
32'h000003af:s1out=32'hcee4c6e8;

32'h000003b0:s1out=32'hef20cada;
32'h000003b1:s1out=32'h36774c01;
32'h000003b2:s1out=32'hd07e9efe;
32'h000003b3:s1out=32'h2bf11fb4;
32'h000003b4:s1out=32'h95dbda4d;
32'h000003b5:s1out=32'hae909198;
32'h000003b6:s1out=32'heaad8e71;
32'h000003b7:s1out=32'h6b93d5a0;
32'h000003b8:s1out=32'hd08ed1d0;
32'h000003b9:s1out=32'hafc725e0;
32'h000003ba:s1out=32'h8e3c5b2f;
32'h000003bb:s1out=32'h8e7594b7;
32'h000003bc:s1out=32'h8ff6e2fb;
32'h000003bd:s1out=32'hf2122b64;
32'h000003be:s1out=32'h8888b812;
32'h000003bf:s1out=32'h900df01c;

32'h000003c0:s1out=32'h4fad5ea0;
32'h000003c1:s1out=32'h688fc32c;
32'h000003c2:s1out=32'hd1cff191;
32'h000003c3:s1out=32'hb3a8c1ad;
32'h000003c4:s1out=32'h2f2f2218;
32'h000003c5:s1out=32'hbe0e1777;
32'h000003c6:s1out=32'hea752dfe;
32'h000003c7:s1out=32'h8b021fa1;
32'h000003c8:s1out=32'he5a0cc0f;
32'h000003c9:s1out=32'hb56f74e8;
32'h000003ca:s1out=32'h18acf3d6;
32'h000003cb:s1out=32'hce89e299;
32'h000003cc:s1out=32'hb4a84fe0;
32'h000003cd:s1out=32'hfd13e0b7;
32'h000003ce:s1out=32'h7cc43b81;
32'h000003cf:s1out=32'hd2ada8d9;

32'h000003d0:s1out=32'h165fa266;
32'h000003d1:s1out=32'h80957705;
32'h000003d2:s1out=32'h93cc7324;
32'h000003d3:s1out=32'h211a1477;
32'h000003d4:s1out=32'he6ad2065;
32'h000003d5:s1out=32'h77b5fa86;
32'h000003d6:s1out=32'hc75442f5;
32'h000003d7:s1out=32'hfb9d35cf;
32'h000003d8:s1out=32'hebcdaf0c;
32'h000003d9:s1out=32'h7b3e89a0;
32'h000003da:s1out=32'hd6411bd3;
32'h000003db:s1out=32'hae1e7e49;
32'h000003dc:s1out=32'h00250e2d;
32'h000003dd:s1out=32'h2071b35e;
32'h000003de:s1out=32'h226800bb;
32'h000003df:s1out=32'h57b8e0af;

32'h000003e0:s1out=32'h2464369b;
32'h000003e1:s1out=32'hf009b91e;
32'h000003e2:s1out=32'h5563911d;
32'h000003e3:s1out=32'h59dfa6aa;
32'h000003e4:s1out=32'h78c14389;
32'h000003e5:s1out=32'hd95a537f;
32'h000003e6:s1out=32'h207d5ba2;
32'h000003e7:s1out=32'h02e5b9c5;
32'h000003e8:s1out=32'h83260376;
32'h000003e9:s1out=32'h6295cfa9;
32'h000003ea:s1out=32'h11c81968;
32'h000003eb:s1out=32'h4e734a41;
32'h000003ec:s1out=32'hb3472dca;
32'h000003ed:s1out=32'h7b14a94a;
32'h000003ee:s1out=32'h1b510052;
32'h000003ef:s1out=32'h9a532915;

32'h000003f0:s1out=32'hd60f573f;
32'h000003f1:s1out=32'hbc9bc6e4;
32'h000003f2:s1out=32'h2b60a476;
32'h000003f3:s1out=32'h81e67400;
32'h000003f4:s1out=32'h08ba6fb5;
32'h000003f5:s1out=32'h571be91f;
32'h000003f6:s1out=32'hf296ec6b;
32'h000003f7:s1out=32'h2a0dd915;
32'h000003f8:s1out=32'hb6636521;
32'h000003f9:s1out=32'he7b9f9b6;
32'h000003fa:s1out=32'hff34052e;
32'h000003fb:s1out=32'hc5855664;
32'h0000003fc:s1out=32'h53b02d5d;
32'h0000003fd:s1out=32'ha99f8fa1;
32'h0000003fe:s1out=32'h08ba4799;
32'h0000003ff:s1out=32'h6e85076a;
 
default:s1out=32'h0000000000; 
endcase
end
pipo_register p1(s1out,clk,rst,sr1out);


endmodule


